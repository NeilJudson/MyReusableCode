library verilog;
use verilog.vl_types.all;
entity multiplier_35 is
    port(
        i_clk           : in     vl_logic;
        i_rst           : in     vl_logic;
        i_en            : in     vl_logic;
        i_a             : in     vl_logic_vector(34 downto 0);
        i_b             : in     vl_logic_vector(34 downto 0);
        o_in_en         : out    vl_logic;
        o_c             : out    vl_logic_vector(68 downto 0);
        o_c_en          : out    vl_logic
    );
end multiplier_35;
